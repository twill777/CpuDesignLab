library verilog;
use verilog.vl_types.all;
entity \Bus\ is
    port(
        BusMuxR0In      : in     vl_logic_vector(31 downto 0);
        BusMuxR1In      : in     vl_logic_vector(31 downto 0);
        BusMuxR2In      : in     vl_logic_vector(31 downto 0);
        BusMuxR3In      : in     vl_logic_vector(31 downto 0);
        BusMuxR4In      : in     vl_logic_vector(31 downto 0);
        BusMuxR5In      : in     vl_logic_vector(31 downto 0);
        BusMuxR6In      : in     vl_logic_vector(31 downto 0);
        BusMuxR7In      : in     vl_logic_vector(31 downto 0);
        BusMuxR8In      : in     vl_logic_vector(31 downto 0);
        BusMuxR9In      : in     vl_logic_vector(31 downto 0);
        BusMuxR10In     : in     vl_logic_vector(31 downto 0);
        BusMuxR11In     : in     vl_logic_vector(31 downto 0);
        BusMuxR12In     : in     vl_logic_vector(31 downto 0);
        BusMuxR13In     : in     vl_logic_vector(31 downto 0);
        BusMuxR14In     : in     vl_logic_vector(31 downto 0);
        BusMuxR15In     : in     vl_logic_vector(31 downto 0);
        BusMuxHIIn      : in     vl_logic_vector(31 downto 0);
        BusMuxLOIn      : in     vl_logic_vector(31 downto 0);
        BusMuxZhighIn   : in     vl_logic_vector(31 downto 0);
        BusMuxZlowIn    : in     vl_logic_vector(31 downto 0);
        BusMuxPCIn      : in     vl_logic_vector(31 downto 0);
        BusMuxMDRIn     : in     vl_logic_vector(31 downto 0);
        BusMuxPortIn    : in     vl_logic_vector(31 downto 0);
        C_sign_extended : in     vl_logic_vector(31 downto 0);
        R0out           : in     vl_logic;
        R1out           : in     vl_logic;
        R2out           : in     vl_logic;
        R3out           : in     vl_logic;
        R4out           : in     vl_logic;
        R5out           : in     vl_logic;
        R6out           : in     vl_logic;
        R7out           : in     vl_logic;
        R8out           : in     vl_logic;
        R9out           : in     vl_logic;
        R10out          : in     vl_logic;
        R11out          : in     vl_logic;
        R12out          : in     vl_logic;
        R13out          : in     vl_logic;
        R14out          : in     vl_logic;
        R15out          : in     vl_logic;
        HIout           : in     vl_logic;
        LOout           : in     vl_logic;
        Zhighout        : in     vl_logic;
        Zlowout         : in     vl_logic;
        PCout           : in     vl_logic;
        MDRout          : in     vl_logic;
        Portout         : in     vl_logic;
        Cout            : in     vl_logic;
        clk             : in     vl_logic;
        BusMuxOut       : out    vl_logic_vector(31 downto 0)
    );
end \Bus\;

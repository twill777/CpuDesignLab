library verilog;
use verilog.vl_types.all;
entity Registers_tb is
end Registers_tb;
